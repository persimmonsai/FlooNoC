

module snitch_cluster_wrapper_test;